LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MAR IS
PORT(
	ADDR_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0); --PCOUT
   IMAR: IN STD_LOGIC;
   CLK: IN STD_LOGIC;
   ADDR_OUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END;

ARCHITECTURE A OF MAR IS
BEGIN 
  PROCESS(CLK,IMAR)
  BEGIN
	IF(CLK'EVENT AND CLK='1') THEN
		IF (IMAR='0') THEN
			ADDR_OUT <= ADDR_IN;
		END IF;
	END IF;
  END PROCESS;
END A;
