library verilog;
use verilog.vl_types.all;
entity CLK_SOURCE_vlg_check_tst is
    port(
        CLK             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CLK_SOURCE_vlg_check_tst;
