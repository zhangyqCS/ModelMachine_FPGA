LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--存储器模块
--可以实现读写功能

ENTITY RAM IS
PORT(
	WR,CS: IN STD_LOGIC;  --CS为片选端，WR为读写端
   DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入指令码
   DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --输出的指令码
   ADDR: IN STD_LOGIC_VECTOR(2 DOWNTO 0) --输入的地址码
);
END;

ARCHITECTURE A OF RAM IS
TYPE MEMORY IS ARRAY(0 TO 4) OF STD_LOGIC_VECTOR(7 DOWNTO 0); --MEMORY为大小为5的数组
BEGIN
   PROCESS(CS,WR)
   VARIABLE MEM:MEMORY;
   BEGIN
      IF(CS='0') THEN
        IF(WR='0') THEN --WR=0进行写入操作
          MEM(CONV_INTEGER(ADDR(2 DOWNTO 0))):=DIN; --强制类型转换为整数
        ELSIF(WR='1') THEN --WR=1进行读出操作
          DOUT <= MEM(CONV_INTEGER(ADDR(2 DOWNTO 0)));
		  END IF;
		END IF;
	END PROCESS;
END A;
