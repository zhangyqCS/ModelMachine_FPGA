library verilog;
use verilog.vl_types.all;
entity COUNTER_vlg_vec_tst is
end COUNTER_vlg_vec_tst;
