library verilog;
use verilog.vl_types.all;
entity Mytest_vlg_vec_tst is
end Mytest_vlg_vec_tst;
