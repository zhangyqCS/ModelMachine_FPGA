library verilog;
use verilog.vl_types.all;
entity ACC_vlg_check_tst is
    port(
        DATA_OUT        : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end ACC_vlg_check_tst;
