library verilog;
use verilog.vl_types.all;
entity COUNTER_vlg_check_tst is
    port(
        T0              : in     vl_logic;
        T1              : in     vl_logic;
        T2              : in     vl_logic;
        T3              : in     vl_logic;
        T4              : in     vl_logic;
        T5              : in     vl_logic;
        T6              : in     vl_logic;
        T7              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end COUNTER_vlg_check_tst;
