library verilog;
use verilog.vl_types.all;
entity RAM_MUX_vlg_vec_tst is
end RAM_MUX_vlg_vec_tst;
