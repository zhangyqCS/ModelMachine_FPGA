library verilog;
use verilog.vl_types.all;
entity MAR_vlg_vec_tst is
end MAR_vlg_vec_tst;
