LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU IS
PORT(
	AC,DR:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	ISUM: IN STD_LOGIC;
	ESUM: IN STD_LOGIC;
	ALU_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END ALU;

ARCHITECTURE A OF ALU IS
SIGNAL ALU_TEMP: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	ALU_TEMP <= AC+DR WHEN ISUM='0';
	ALU_OUT <= ALU_TEMP WHEN ESUM='0';
	
	--ALU_OUT <= CONV_INTEGER(ALU_TEMP(7 DOWNTO 0));
END A;
