LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--数据选择器
--可以实现手动向存储器制定地址单元写入数据

ENTITY RAM_MUX IS
PORT(
	SEL : IN STD_LOGIC;
	DATA0X : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	DATA1X : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	RESULT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);

END;

ARCHITECTURE A OF RAM_MUX IS
BEGIN

	RESULT <= DATA0X WHEN SEL='0' ELSE DATA1X; 
	
END A;
	