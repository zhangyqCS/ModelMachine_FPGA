library verilog;
use verilog.vl_types.all;
entity ACC_vlg_vec_tst is
end ACC_vlg_vec_tst;
