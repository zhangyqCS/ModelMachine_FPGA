library verilog;
use verilog.vl_types.all;
entity RAM_vlg_vec_tst is
end RAM_vlg_vec_tst;
