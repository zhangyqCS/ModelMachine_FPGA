LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

--地址寄存器模块
--临时存放地址码

ENTITY MAR IS
PORT(
	ADDR_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0); --从PC接收的地址码
   IMAR: IN STD_LOGIC; --MAR允许输出信号
   CLK: IN STD_LOGIC; --时钟信号
   ADDR_OUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0) --MAR输出地址码端口
);
END;

ARCHITECTURE A OF MAR IS
BEGIN 
  PROCESS(CLK,IMAR)
  BEGIN
	IF(CLK'EVENT AND CLK='1') THEN --CLK上升沿到来时
		IF (IMAR='0') THEN  --IMAR=0时允许输出
			ADDR_OUT <= ADDR_IN;
		END IF;
	END IF;
  END PROCESS;
END A;
