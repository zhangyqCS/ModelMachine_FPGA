library verilog;
use verilog.vl_types.all;
entity DR_vlg_vec_tst is
end DR_vlg_vec_tst;
