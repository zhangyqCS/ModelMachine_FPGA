library verilog;
use verilog.vl_types.all;
entity MC_TEMP_vlg_vec_tst is
end MC_TEMP_vlg_vec_tst;
