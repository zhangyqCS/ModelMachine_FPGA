LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RAM IS
PORT(
	--WR,CS: IN STD_LOGIC;
   --DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
   DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
   ADDR: IN STD_LOGIC_VECTOR(2 DOWNTO 0) --MAR_OUT
);
END;

ARCHITECTURE A OF RAM IS
TYPE MEMORY IS ARRAY(0 TO 4) OF STD_LOGIC_VECTOR(7 DOWNTO 0); --MEMORY为数组
--SIGNAL MEMY : MEMORY;
--VARIABLE MEM:MEMORY;
BEGIN
	--MEM(0) := "00111110";
	--MEM(1) := "00000110";
	--MEM(2) := "11000110";
	--MEM(3) := "00000111";
	--MEM(4) := "01110110";
   PROCESS(ADDR)
   VARIABLE MEM:MEMORY;
   BEGIN
	MEM(0) := "00111110";
	MEM(1) := "00000010";
	MEM(2) := "11000110";
	MEM(3) := "00000111";
	MEM(4) := "01110110";
      --IF(CS='0') THEN
        --IF(WR='0') THEN
          --MEM(CONV_INTEGER(ADDR(2 DOWNTO 0))) :=DIN; --强制类型转换为整数
        --IF(WR='1') THEN
          DOUT <= MEM(CONV_INTEGER(ADDR(2 DOWNTO 0)));
		  --END IF;
		--END IF;
	END PROCESS;
END A;
