library verilog;
use verilog.vl_types.all;
entity IR_vlg_vec_tst is
end IR_vlg_vec_tst;
