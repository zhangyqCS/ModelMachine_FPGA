LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--算数逻辑单元
--可以实现两个立即数相加并将结果输出

ENTITY ALU IS
PORT(
	AC,DR:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入的两个立即数
	ISUM: IN STD_LOGIC; --ALU加法操作信号
	ESUM: IN STD_LOGIC; --ALU允许输出信号
	ALU_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0) --输出结果信号
);
END ALU;

ARCHITECTURE A OF ALU IS
SIGNAL ALU_TEMP: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	ALU_TEMP <= AC+DR WHEN ISUM='0'; --ISUM=0时实现两个立即数相加
	ALU_OUT <= ALU_TEMP WHEN ESUM='0'; --ESUM=0输出。
END A;
