LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--程序计数器模块
--用以产生正确的地址

ENTITY PC IS
PORT( 
	IPC,CLK,CLR: IN STD_LOGIC; --CLK为时钟周期，CLR为复位端，IPC为允许计数指令
   PCOUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0) --输出产生的地址码
);
END;

ARCHITECTURE A OF PC IS
SIGNAL QOUT: STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN
PROCESS(CLK,CLR,IPC)
BEGIN
   IF(CLR='0') THEN  --CLR=0时复位，将000赋值给QOUT
      QOUT <= "000";
   ELSIF(CLK'EVENT AND CLK='1') THEN --CLK上升沿
      IF(IPC='1') THEN --IPC=1时程序计数
			QOUT <= QOUT+1; --QOUT执行QOUT+1操作
      END IF;
   END IF;
END PROCESS;
  PCOUT<=QOUT;
END A;
