LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PC IS
PORT( 
	IPC,CLK,CLR: IN STD_LOGIC;
   PCOUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END;

ARCHITECTURE A OF PC IS
SIGNAL QOUT: STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN
PROCESS(CLK,CLR,IPC)
BEGIN
   IF(CLR='0') THEN
      QOUT <= "000";
   ELSIF(CLK'EVENT AND CLK='1') THEN
      IF(IPC='1') THEN
			QOUT <= QOUT+1;
      END IF;
   END IF;
END PROCESS;
  PCOUT<=QOUT;
END A;
