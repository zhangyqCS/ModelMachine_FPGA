library verilog;
use verilog.vl_types.all;
entity CLK_SOURCE_vlg_vec_tst is
end CLK_SOURCE_vlg_vec_tst;
