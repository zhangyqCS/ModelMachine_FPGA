library verilog;
use verilog.vl_types.all;
entity CTRL_vlg_vec_tst is
end CTRL_vlg_vec_tst;
