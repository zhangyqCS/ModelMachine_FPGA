library verilog;
use verilog.vl_types.all;
entity DR_vlg_check_tst is
    port(
        DATA_OUT        : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end DR_vlg_check_tst;
